
module preamble_detect # (
    parameter SAMPLE_RATE = 16,
    parameter TRANSITION_ERROR = 1
) (
    input logic clk,
    input logic en,
    input logic resetn,

    input logic data_bit,
    output logic preamble_detected
);

    localparam PREAMBLE_LEN = 8;
    localparam BUFFER_LEN = (PREAMBLE_LEN - 1) * SAMPLE_RATE + 2 * TRANSITION_ERROR - 1;
    // Buffer to store when matched filter output transitions occur in the last (PREAMBLE_LEN-1) * SAMPLE_RATE + TRANSITION_ERROR - 1 cycles
    logic [BUFFER_LEN-1:0] transition_buffer;
    logic last_bit, valid_transition;
    int i, j;

    always_comb begin
        // A preamble is detected if the matched filter output transitions on the current clock cycle and within TRANSITION_ERROR sample(s) of the previous cycles where CYCLE % SAMPLE_RATE == SAMPLE_RATE - 1
        preamble_detected = data_bit ^ last_bit;
        for (i = SAMPLE_RATE - 1; i < BUFFER_LEN; i = i + SAMPLE_RATE) begin
            valid_transition = 1'b0;
            for (j = -TRANSITION_ERROR; j <= TRANSITION_ERROR; j = j + 1) begin
                valid_transition = valid_transition ^ transition_buffer[i + j];
            end

            preamble_detected = preamble_detected & valid_transition;
        end
    end

    always_ff @(posedge clk or negedge resetn) begin
        if (~resetn) begin
            transition_buffer <= {BUFFER_LEN{1'b0}};
            last_bit <= 0;
        end else if (en) begin
            // Shift the buffer, and store if the matched filter output transitions. Keep track of the previous bit
            transition_buffer <= {transition_buffer[BUFFER_LEN-2:0], data_bit ^ last_bit};
            last_bit <= data_bit;
        end
    end

endmodule

